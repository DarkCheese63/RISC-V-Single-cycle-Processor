-------------------------------------------------------------------------
-- Matthew Estes
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------
-- tb_ALUControl.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: this is the test bench for the ALU control
--              
-- 10/21/2025
-------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb_ALUControl is
end tb_ALUControl;




